module SB_SPRAM256KA(
	ADDRESS, DATAIN, MASKWREN,WREN,CHIPSELECT,CLOCK,STANDBY,SLEEP,POWEROFF,DATAOUT
)/* synthesis syn_black_box syn_lib_cell=1 TEST_SPRAM="" */;
input [13:0] ADDRESS;
input [15:0] DATAIN;
input [3:0] MASKWREN;
input WREN,CHIPSELECT,CLOCK,STANDBY,SLEEP,POWEROFF;
output [15:0] DATAOUT;
endmodule
 