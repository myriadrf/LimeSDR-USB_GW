@00000000
18000000
18400000
18A00000
18200000
A8210000
BC010000
0FFFFFFF
9C21FFFF
1880B000
A8400051
D8041000
D8040004
A8C00001
D8043004
A8A00001
04000022
A8600003
04000020
A8600000
0400001E
A8600000
0400001C
A860000C
A8A00004
04000019
15000000
E1620004
04000016
15000000
E1820004
04000013
15000000
E1A20004
A8C00009
0400000F
15000000
BC060000
0FFFFFFD
9CC6FFFF
18C00000
04000009
E0EC3000
D4071000
9CC60004
E4665800
0FFFFFFB
15000000
44006800
D8040004
E0250004
D8041802
A8600001
A4630001
BC030001
13FFFFFE
8C640001
8C640002
B8420008
E0421804
BC010001
0FFFFFF6
9C21FFFF
44004800
15000000
