-- lms_orca.vhd

-- Generated using ACDS version 15.1 193

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lms_orca is
	port (
		clk_clk                                     : in    std_logic                     := '0';             --                                  clk.clk
		controlled_reset_external_connection_export : out   std_logic;                                        -- controlled_reset_external_connection.export
		exfifo_if_d_export                          : in    std_logic_vector(31 downto 0) := (others => '0'); --                          exfifo_if_d.export
		exfifo_if_rd_export                         : out   std_logic;                                        --                         exfifo_if_rd.export
		exfifo_if_rdempty_export                    : in    std_logic                     := '0';             --                    exfifo_if_rdempty.export
		exfifo_of_d_export                          : out   std_logic_vector(31 downto 0);                    --                          exfifo_of_d.export
		exfifo_of_wr_export                         : out   std_logic;                                        --                         exfifo_of_wr.export
		exfifo_of_wrfull_export                     : in    std_logic                     := '0';             --                     exfifo_of_wrfull.export
		exfifo_rst_export                           : out   std_logic;                                        --                           exfifo_rst.export
		i2c_opencores_0_interrupt_sender_irq        : out   std_logic;                                        --     i2c_opencores_0_interrupt_sender.irq
		in_reset_reset_n                            : in    std_logic                     := '0';             --                             in_reset.reset_n
		leds_external_connection_export             : out   std_logic_vector(7 downto 0);                     --             leds_external_connection.export
		lms_ctr_gpio_external_connection_export     : out   std_logic_vector(3 downto 0);                     --     lms_ctr_gpio_external_connection.export
		scl_exp_export                              : inout std_logic                     := '0';             --                              scl_exp.export
		sda_exp_export                              : inout std_logic                     := '0';             --                              sda_exp.export
		spi_1_dac_external_MISO                     : in    std_logic                     := '0';             --                   spi_1_dac_external.MISO
		spi_1_dac_external_MOSI                     : out   std_logic;                                        --                                     .MOSI
		spi_1_dac_external_SCLK                     : out   std_logic;                                        --                                     .SCLK
		spi_1_dac_external_SS_n                     : out   std_logic_vector(1 downto 0);                     --                                     .SS_n
		spi_1_dac_irq_irq                           : out   std_logic;                                        --                        spi_1_dac_irq.irq
		spi_lms_external_MISO                       : in    std_logic                     := '0';             --                     spi_lms_external.MISO
		spi_lms_external_MOSI                       : out   std_logic;                                        --                                     .MOSI
		spi_lms_external_SCLK                       : out   std_logic;                                        --                                     .SCLK
		spi_lms_external_SS_n                       : out   std_logic_vector(4 downto 0);                     --                                     .SS_n
		spi_lms_irq_irq                             : out   std_logic;                                        --                          spi_lms_irq.irq
		switch_external_connection_export           : in    std_logic_vector(7 downto 0)  := (others => '0'); --           switch_external_connection.export
		vectorblox_orca_0_global_interrupts_export  : in    std_logic_vector(0 downto 0)  := (others => '0')  --  vectorblox_orca_0_global_interrupts.export
	);
end entity lms_orca;

architecture rtl of lms_orca is
	component avfifo is
		generic (
			width : integer := 32
		);
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect     : in  std_logic                     := 'X';             -- chipselect
			write          : in  std_logic                     := 'X';             -- write
			writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read           : in  std_logic                     := 'X';             -- read
			readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			rsi_nrst       : in  std_logic                     := 'X';             -- reset_n
			coe_if_d       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			coe_if_rd      : out std_logic;                                        -- export
			coe_of_wrfull  : in  std_logic                     := 'X';             -- export
			coe_of_wr      : out std_logic;                                        -- export
			coe_of_d       : out std_logic_vector(31 downto 0);                    -- export
			coe_if_rdempty : in  std_logic                     := 'X';             -- export
			coe_fifo_rst   : out std_logic                                         -- export
		);
	end component avfifo;

	component lms_orca_controlled_reset is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component lms_orca_controlled_reset;

	component i2c_opencores is
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component i2c_opencores;

	component lms_orca_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component lms_orca_leds;

	component lms_orca_lms_ctr_gpio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component lms_orca_lms_ctr_gpio;

	component lms_orca_oc_mem is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component lms_orca_oc_mem;

	component lms_orca_spi_1_DAC is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic_vector(1 downto 0)                      -- export
		);
	end component lms_orca_spi_1_DAC;

	component lms_orca_spi_lms is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic_vector(4 downto 0)                      -- export
		);
	end component lms_orca_spi_lms;

	component lms_orca_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component lms_orca_switch;

	component lms_orca_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component lms_orca_sysid_qsys_0;

	component Orca is
		generic (
			REGISTER_SIZE         : integer := 32;
			AVALON_ENABLE         : natural := 1;
			AXI_ENABLE            : natural := 0;
			LVE_ENABLE            : natural := 0;
			SCRATCHPAD_SIZE       : integer := 1024;
			RESET_VECTOR          : integer := 512;
			MULTIPLY_ENABLE       : natural := 0;
			DIVIDE_ENABLE         : natural := 0;
			SHIFTER_MAX_CYCLES    : natural := 32;
			ENABLE_EXCEPTIONS     : natural := 1;
			NUM_EXT_INTERRUPTS    : integer := 1;
			ENABLE_EXT_INTERRUPTS : natural := 1;
			COUNTER_LENGTH        : natural := 64;
			BRANCH_PREDICTORS     : natural := 1;
			PIPELINE_STAGES       : natural := 4
		);
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			scratchpad_clk                : in  std_logic                     := 'X';             -- clk
			reset                         : in  std_logic                     := 'X';             -- reset
			avm_data_address              : out std_logic_vector(31 downto 0);                    -- address
			avm_data_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_data_read                 : out std_logic;                                        -- read
			avm_data_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_data_write                : out std_logic;                                        -- write
			avm_data_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			avm_data_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			avm_data_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			data_ARADDR                   : out std_logic_vector(31 downto 0);                    -- araddr
			data_ARBURST                  : out std_logic_vector(1 downto 0);                     -- arburst
			data_ARCACHE                  : out std_logic_vector(3 downto 0);                     -- arcache
			data_ARID                     : out std_logic_vector(3 downto 0);                     -- arid
			data_ARLEN                    : out std_logic_vector(3 downto 0);                     -- arlen
			data_ARLOCK                   : out std_logic_vector(1 downto 0);                     -- arlock
			data_ARPROT                   : out std_logic_vector(2 downto 0);                     -- arprot
			data_ARREADY                  : in  std_logic                     := 'X';             -- arready
			data_ARSIZE                   : out std_logic_vector(2 downto 0);                     -- arsize
			data_ARVALID                  : out std_logic;                                        -- arvalid
			data_AWADDR                   : out std_logic_vector(31 downto 0);                    -- awaddr
			data_AWBURST                  : out std_logic_vector(1 downto 0);                     -- awburst
			data_AWCACHE                  : out std_logic_vector(3 downto 0);                     -- awcache
			data_AWID                     : out std_logic_vector(3 downto 0);                     -- awid
			data_AWLEN                    : out std_logic_vector(3 downto 0);                     -- awlen
			data_AWLOCK                   : out std_logic_vector(1 downto 0);                     -- awlock
			data_AWPROT                   : out std_logic_vector(2 downto 0);                     -- awprot
			data_AWREADY                  : in  std_logic                     := 'X';             -- awready
			data_AWSIZE                   : out std_logic_vector(2 downto 0);                     -- awsize
			data_AWVALID                  : out std_logic;                                        -- awvalid
			data_BID                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- bid
			data_BREADY                   : out std_logic;                                        -- bready
			data_BRESP                    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			data_BVALID                   : in  std_logic                     := 'X';             -- bvalid
			data_RDATA                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			data_RID                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rid
			data_RLAST                    : in  std_logic                     := 'X';             -- rlast
			data_RREADY                   : out std_logic;                                        -- rready
			data_RRESP                    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			data_RVALID                   : in  std_logic                     := 'X';             -- rvalid
			data_WDATA                    : out std_logic_vector(31 downto 0);                    -- wdata
			data_WID                      : out std_logic_vector(3 downto 0);                     -- wid
			data_WLAST                    : out std_logic;                                        -- wlast
			data_WREADY                   : in  std_logic                     := 'X';             -- wready
			data_WSTRB                    : out std_logic_vector(3 downto 0);                     -- wstrb
			data_WVALID                   : out std_logic;                                        -- wvalid
			instr_ARADDR                  : out std_logic_vector(31 downto 0);                    -- araddr
			instr_ARBURST                 : out std_logic_vector(1 downto 0);                     -- arburst
			instr_ARCACHE                 : out std_logic_vector(3 downto 0);                     -- arcache
			instr_ARID                    : out std_logic_vector(3 downto 0);                     -- arid
			instr_ARLEN                   : out std_logic_vector(3 downto 0);                     -- arlen
			instr_ARLOCK                  : out std_logic_vector(1 downto 0);                     -- arlock
			instr_ARPROT                  : out std_logic_vector(2 downto 0);                     -- arprot
			instr_ARREADY                 : in  std_logic                     := 'X';             -- arready
			instr_ARSIZE                  : out std_logic_vector(2 downto 0);                     -- arsize
			instr_ARVALID                 : out std_logic;                                        -- arvalid
			instr_AWADDR                  : out std_logic_vector(31 downto 0);                    -- awaddr
			instr_AWBURST                 : out std_logic_vector(1 downto 0);                     -- awburst
			instr_AWCACHE                 : out std_logic_vector(3 downto 0);                     -- awcache
			instr_AWID                    : out std_logic_vector(3 downto 0);                     -- awid
			instr_AWLEN                   : out std_logic_vector(3 downto 0);                     -- awlen
			instr_AWLOCK                  : out std_logic_vector(1 downto 0);                     -- awlock
			instr_AWPROT                  : out std_logic_vector(2 downto 0);                     -- awprot
			instr_AWREADY                 : in  std_logic                     := 'X';             -- awready
			instr_AWSIZE                  : out std_logic_vector(2 downto 0);                     -- awsize
			instr_AWVALID                 : out std_logic;                                        -- awvalid
			instr_BID                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- bid
			instr_BREADY                  : out std_logic;                                        -- bready
			instr_BRESP                   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			instr_BVALID                  : in  std_logic                     := 'X';             -- bvalid
			instr_RDATA                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			instr_RID                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rid
			instr_RLAST                   : in  std_logic                     := 'X';             -- rlast
			instr_RREADY                  : out std_logic;                                        -- rready
			instr_RRESP                   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			instr_RVALID                  : in  std_logic                     := 'X';             -- rvalid
			instr_WDATA                   : out std_logic_vector(31 downto 0);                    -- wdata
			instr_WID                     : out std_logic_vector(3 downto 0);                     -- wid
			instr_WLAST                   : out std_logic;                                        -- wlast
			instr_WREADY                  : in  std_logic                     := 'X';             -- wready
			instr_WSTRB                   : out std_logic_vector(3 downto 0);                     -- wstrb
			instr_WVALID                  : out std_logic;                                        -- wvalid
			avm_instruction_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_instruction_read          : out std_logic;                                        -- read
			avm_instruction_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_instruction_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_instruction_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			global_interrupts             : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- export
			data_ADR_O                    : out std_logic_vector(31 downto 0);                    -- export0
			data_DAT_I                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export1
			data_DAT_O                    : out std_logic_vector(31 downto 0);                    -- export2
			data_WE_O                     : out std_logic;                                        -- export3
			data_SEL_O                    : out std_logic_vector(3 downto 0);                     -- export4
			data_STB_O                    : out std_logic;                                        -- export5
			data_ACK_I                    : in  std_logic                     := 'X';             -- export6
			data_CYC_O                    : out std_logic;                                        -- export7
			data_CTI_O                    : out std_logic_vector(2 downto 0);                     -- export8
			data_STALL_I                  : in  std_logic                     := 'X';             -- export9
			instr_ADR_O                   : out std_logic_vector(31 downto 0);                    -- export10
			instr_DAT_I                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export11
			instr_STB_O                   : out std_logic;                                        -- export12
			instr_ACK_I                   : in  std_logic                     := 'X';             -- export13
			instr_CYC_O                   : out std_logic;                                        -- export14
			instr_CTI_O                   : out std_logic_vector(2 downto 0);                     -- export15
			instr_STALL_I                 : in  std_logic                     := 'X'              -- export16
		);
	end component Orca;

	component lms_orca_mm_interconnect_0 is
		port (
			clk_main_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			vectorblox_orca_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			vectorblox_orca_0_data_address                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vectorblox_orca_0_data_waitrequest                  : out std_logic;                                        -- waitrequest
			vectorblox_orca_0_data_byteenable                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			vectorblox_orca_0_data_read                         : in  std_logic                     := 'X';             -- read
			vectorblox_orca_0_data_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			vectorblox_orca_0_data_readdatavalid                : out std_logic;                                        -- readdatavalid
			vectorblox_orca_0_data_write                        : in  std_logic                     := 'X';             -- write
			vectorblox_orca_0_data_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			vectorblox_orca_0_instruction_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vectorblox_orca_0_instruction_waitrequest           : out std_logic;                                        -- waitrequest
			vectorblox_orca_0_instruction_read                  : in  std_logic                     := 'X';             -- read
			vectorblox_orca_0_instruction_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			vectorblox_orca_0_instruction_readdatavalid         : out std_logic;                                        -- readdatavalid
			Av_FIFO_Int_0_avalon_slave_0_address                : out std_logic_vector(1 downto 0);                     -- address
			Av_FIFO_Int_0_avalon_slave_0_write                  : out std_logic;                                        -- write
			Av_FIFO_Int_0_avalon_slave_0_read                   : out std_logic;                                        -- read
			Av_FIFO_Int_0_avalon_slave_0_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Av_FIFO_Int_0_avalon_slave_0_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			Av_FIFO_Int_0_avalon_slave_0_chipselect             : out std_logic;                                        -- chipselect
			controlled_reset_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			controlled_reset_s1_write                           : out std_logic;                                        -- write
			controlled_reset_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			controlled_reset_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			controlled_reset_s1_chipselect                      : out std_logic;                                        -- chipselect
			i2c_opencores_0_avalon_slave_0_address              : out std_logic_vector(2 downto 0);                     -- address
			i2c_opencores_0_avalon_slave_0_write                : out std_logic;                                        -- write
			i2c_opencores_0_avalon_slave_0_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_opencores_0_avalon_slave_0_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_opencores_0_avalon_slave_0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect           : out std_logic;                                        -- chipselect
			leds_s1_address                                     : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                       : out std_logic;                                        -- write
			leds_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                                  : out std_logic;                                        -- chipselect
			lms_ctr_gpio_s1_address                             : out std_logic_vector(2 downto 0);                     -- address
			lms_ctr_gpio_s1_write                               : out std_logic;                                        -- write
			lms_ctr_gpio_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lms_ctr_gpio_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			lms_ctr_gpio_s1_chipselect                          : out std_logic;                                        -- chipselect
			oc_mem_s1_address                                   : out std_logic_vector(12 downto 0);                    -- address
			oc_mem_s1_write                                     : out std_logic;                                        -- write
			oc_mem_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			oc_mem_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			oc_mem_s1_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			oc_mem_s1_chipselect                                : out std_logic;                                        -- chipselect
			oc_mem_s1_clken                                     : out std_logic;                                        -- clken
			spi_1_DAC_spi_control_port_address                  : out std_logic_vector(2 downto 0);                     -- address
			spi_1_DAC_spi_control_port_write                    : out std_logic;                                        -- write
			spi_1_DAC_spi_control_port_read                     : out std_logic;                                        -- read
			spi_1_DAC_spi_control_port_readdata                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_1_DAC_spi_control_port_writedata                : out std_logic_vector(15 downto 0);                    -- writedata
			spi_1_DAC_spi_control_port_chipselect               : out std_logic;                                        -- chipselect
			spi_lms_spi_control_port_address                    : out std_logic_vector(2 downto 0);                     -- address
			spi_lms_spi_control_port_write                      : out std_logic;                                        -- write
			spi_lms_spi_control_port_read                       : out std_logic;                                        -- read
			spi_lms_spi_control_port_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_lms_spi_control_port_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			spi_lms_spi_control_port_chipselect                 : out std_logic;                                        -- chipselect
			switch_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_0_control_slave_address                  : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component lms_orca_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal vectorblox_orca_0_data_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:vectorblox_orca_0_data_readdata -> vectorblox_orca_0:avm_data_readdata
	signal vectorblox_orca_0_data_waitrequest                           : std_logic;                     -- mm_interconnect_0:vectorblox_orca_0_data_waitrequest -> vectorblox_orca_0:avm_data_waitrequest
	signal vectorblox_orca_0_data_address                               : std_logic_vector(31 downto 0); -- vectorblox_orca_0:avm_data_address -> mm_interconnect_0:vectorblox_orca_0_data_address
	signal vectorblox_orca_0_data_byteenable                            : std_logic_vector(3 downto 0);  -- vectorblox_orca_0:avm_data_byteenable -> mm_interconnect_0:vectorblox_orca_0_data_byteenable
	signal vectorblox_orca_0_data_read                                  : std_logic;                     -- vectorblox_orca_0:avm_data_read -> mm_interconnect_0:vectorblox_orca_0_data_read
	signal vectorblox_orca_0_data_readdatavalid                         : std_logic;                     -- mm_interconnect_0:vectorblox_orca_0_data_readdatavalid -> vectorblox_orca_0:avm_data_readdatavalid
	signal vectorblox_orca_0_data_write                                 : std_logic;                     -- vectorblox_orca_0:avm_data_write -> mm_interconnect_0:vectorblox_orca_0_data_write
	signal vectorblox_orca_0_data_writedata                             : std_logic_vector(31 downto 0); -- vectorblox_orca_0:avm_data_writedata -> mm_interconnect_0:vectorblox_orca_0_data_writedata
	signal vectorblox_orca_0_instruction_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:vectorblox_orca_0_instruction_readdata -> vectorblox_orca_0:avm_instruction_readdata
	signal vectorblox_orca_0_instruction_waitrequest                    : std_logic;                     -- mm_interconnect_0:vectorblox_orca_0_instruction_waitrequest -> vectorblox_orca_0:avm_instruction_waitrequest
	signal vectorblox_orca_0_instruction_address                        : std_logic_vector(31 downto 0); -- vectorblox_orca_0:avm_instruction_address -> mm_interconnect_0:vectorblox_orca_0_instruction_address
	signal vectorblox_orca_0_instruction_read                           : std_logic;                     -- vectorblox_orca_0:avm_instruction_read -> mm_interconnect_0:vectorblox_orca_0_instruction_read
	signal vectorblox_orca_0_instruction_readdatavalid                  : std_logic;                     -- mm_interconnect_0:vectorblox_orca_0_instruction_readdatavalid -> vectorblox_orca_0:avm_instruction_readdatavalid
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect  : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata    : std_logic_vector(7 downto 0);  -- i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	signal i2c_opencores_0_avalon_slave_0_waitrequest                   : std_logic;                     -- i2c_opencores_0:wb_ack_o -> i2c_opencores_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write       : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect    : std_logic;                     -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_chipselect -> Av_FIFO_Int_0:chipselect
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata      : std_logic_vector(31 downto 0); -- Av_FIFO_Int_0:readdata -> mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_readdata
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_address -> Av_FIFO_Int_0:address
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read          : std_logic;                     -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_read -> Av_FIFO_Int_0:read
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write         : std_logic;                     -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_write -> Av_FIFO_Int_0:write
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_writedata -> Av_FIFO_Int_0:writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata        : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_oc_mem_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:oc_mem_s1_chipselect -> oc_mem:chipselect
	signal mm_interconnect_0_oc_mem_s1_readdata                         : std_logic_vector(31 downto 0); -- oc_mem:readdata -> mm_interconnect_0:oc_mem_s1_readdata
	signal mm_interconnect_0_oc_mem_s1_address                          : std_logic_vector(12 downto 0); -- mm_interconnect_0:oc_mem_s1_address -> oc_mem:address
	signal mm_interconnect_0_oc_mem_s1_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:oc_mem_s1_byteenable -> oc_mem:byteenable
	signal mm_interconnect_0_oc_mem_s1_write                            : std_logic;                     -- mm_interconnect_0:oc_mem_s1_write -> oc_mem:write
	signal mm_interconnect_0_oc_mem_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:oc_mem_s1_writedata -> oc_mem:writedata
	signal mm_interconnect_0_oc_mem_s1_clken                            : std_logic;                     -- mm_interconnect_0:oc_mem_s1_clken -> oc_mem:clken
	signal mm_interconnect_0_lms_ctr_gpio_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:lms_ctr_gpio_s1_chipselect -> lms_ctr_gpio:chipselect
	signal mm_interconnect_0_lms_ctr_gpio_s1_readdata                   : std_logic_vector(31 downto 0); -- lms_ctr_gpio:readdata -> mm_interconnect_0:lms_ctr_gpio_s1_readdata
	signal mm_interconnect_0_lms_ctr_gpio_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:lms_ctr_gpio_s1_address -> lms_ctr_gpio:address
	signal mm_interconnect_0_lms_ctr_gpio_s1_write                      : std_logic;                     -- mm_interconnect_0:lms_ctr_gpio_s1_write -> mm_interconnect_0_lms_ctr_gpio_s1_write:in
	signal mm_interconnect_0_lms_ctr_gpio_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:lms_ctr_gpio_s1_writedata -> lms_ctr_gpio:writedata
	signal mm_interconnect_0_leds_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                           : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                              : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_switch_s1_readdata                         : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_controlled_reset_s1_chipselect             : std_logic;                     -- mm_interconnect_0:controlled_reset_s1_chipselect -> controlled_reset:chipselect
	signal mm_interconnect_0_controlled_reset_s1_readdata               : std_logic_vector(31 downto 0); -- controlled_reset:readdata -> mm_interconnect_0:controlled_reset_s1_readdata
	signal mm_interconnect_0_controlled_reset_s1_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:controlled_reset_s1_address -> controlled_reset:address
	signal mm_interconnect_0_controlled_reset_s1_write                  : std_logic;                     -- mm_interconnect_0:controlled_reset_s1_write -> mm_interconnect_0_controlled_reset_s1_write:in
	signal mm_interconnect_0_controlled_reset_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:controlled_reset_s1_writedata -> controlled_reset:writedata
	signal mm_interconnect_0_spi_1_dac_spi_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:spi_1_DAC_spi_control_port_chipselect -> spi_1_DAC:spi_select
	signal mm_interconnect_0_spi_1_dac_spi_control_port_readdata        : std_logic_vector(15 downto 0); -- spi_1_DAC:data_to_cpu -> mm_interconnect_0:spi_1_DAC_spi_control_port_readdata
	signal mm_interconnect_0_spi_1_dac_spi_control_port_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_1_DAC_spi_control_port_address -> spi_1_DAC:mem_addr
	signal mm_interconnect_0_spi_1_dac_spi_control_port_read            : std_logic;                     -- mm_interconnect_0:spi_1_DAC_spi_control_port_read -> mm_interconnect_0_spi_1_dac_spi_control_port_read:in
	signal mm_interconnect_0_spi_1_dac_spi_control_port_write           : std_logic;                     -- mm_interconnect_0:spi_1_DAC_spi_control_port_write -> mm_interconnect_0_spi_1_dac_spi_control_port_write:in
	signal mm_interconnect_0_spi_1_dac_spi_control_port_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_1_DAC_spi_control_port_writedata -> spi_1_DAC:data_from_cpu
	signal mm_interconnect_0_spi_lms_spi_control_port_chipselect        : std_logic;                     -- mm_interconnect_0:spi_lms_spi_control_port_chipselect -> spi_lms:spi_select
	signal mm_interconnect_0_spi_lms_spi_control_port_readdata          : std_logic_vector(15 downto 0); -- spi_lms:data_to_cpu -> mm_interconnect_0:spi_lms_spi_control_port_readdata
	signal mm_interconnect_0_spi_lms_spi_control_port_address           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_lms_spi_control_port_address -> spi_lms:mem_addr
	signal mm_interconnect_0_spi_lms_spi_control_port_read              : std_logic;                     -- mm_interconnect_0:spi_lms_spi_control_port_read -> mm_interconnect_0_spi_lms_spi_control_port_read:in
	signal mm_interconnect_0_spi_lms_spi_control_port_write             : std_logic;                     -- mm_interconnect_0:spi_lms_spi_control_port_write -> mm_interconnect_0_spi_lms_spi_control_port_write:in
	signal mm_interconnect_0_spi_lms_spi_control_port_writedata         : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_lms_spi_control_port_writedata -> spi_lms:data_from_cpu
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [i2c_opencores_0:wb_rst_i, mm_interconnect_0:vectorblox_orca_0_reset_reset_bridge_in_reset_reset, oc_mem:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, vectorblox_orca_0:reset]
	signal rst_controller_reset_out_reset_req                           : std_logic;                     -- rst_controller:reset_req -> [oc_mem:reset_req, rst_translator:reset_req_in]
	signal in_reset_reset_n_ports_inv                                   : std_logic;                     -- in_reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv         : std_logic;                     -- i2c_opencores_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_lms_ctr_gpio_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_lms_ctr_gpio_s1_write:inv -> lms_ctr_gpio:write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_0_controlled_reset_s1_write_ports_inv        : std_logic;                     -- mm_interconnect_0_controlled_reset_s1_write:inv -> controlled_reset:write_n
	signal mm_interconnect_0_spi_1_dac_spi_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_spi_1_dac_spi_control_port_read:inv -> spi_1_DAC:read_n
	signal mm_interconnect_0_spi_1_dac_spi_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_spi_1_dac_spi_control_port_write:inv -> spi_1_DAC:write_n
	signal mm_interconnect_0_spi_lms_spi_control_port_read_ports_inv    : std_logic;                     -- mm_interconnect_0_spi_lms_spi_control_port_read:inv -> spi_lms:read_n
	signal mm_interconnect_0_spi_lms_spi_control_port_write_ports_inv   : std_logic;                     -- mm_interconnect_0_spi_lms_spi_control_port_write:inv -> spi_lms:write_n
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Av_FIFO_Int_0:rsi_nrst, controlled_reset:reset_n, leds:reset_n, lms_ctr_gpio:reset_n, spi_1_DAC:reset_n, spi_lms:reset_n, switch:reset_n, sysid_qsys_0:reset_n]

begin

	av_fifo_int_0 : component avfifo
		generic map (
			width => 32
		)
		port map (
			clk            => clk_clk,                                                   --          clock.clk
			address        => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address,    -- avalon_slave_0.address
			chipselect     => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect, --               .chipselect
			write          => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write,      --               .write
			writedata      => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata,  --               .writedata
			read           => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read,       --               .read
			readdata       => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata,   --               .readdata
			rsi_nrst       => rst_controller_reset_out_reset_ports_inv,                  --          reset.reset_n
			coe_if_d       => exfifo_if_d_export,                                        --       cnd_if_d.export
			coe_if_rd      => exfifo_if_rd_export,                                       --      cnd_if_rd.export
			coe_of_wrfull  => exfifo_of_wrfull_export,                                   --  cnd_of_wrfull.export
			coe_of_wr      => exfifo_of_wr_export,                                       --      cnd_of_wr.export
			coe_of_d       => exfifo_of_d_export,                                        --       cnd_of_d.export
			coe_if_rdempty => exfifo_if_rdempty_export,                                  -- cnd_if_rdempty.export
			coe_fifo_rst   => exfifo_rst_export                                          --   cnd_fifo_rst.export
		);

	controlled_reset : component lms_orca_controlled_reset
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_controlled_reset_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_controlled_reset_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_controlled_reset_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_controlled_reset_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_controlled_reset_s1_readdata,        --                    .readdata
			out_port   => controlled_reset_external_connection_export            -- external_connection.export
		);

	i2c_opencores_0 : component i2c_opencores
		port map (
			wb_clk_i   => clk_clk,                                                     --            clock.clk
			wb_rst_i   => rst_controller_reset_out_reset,                              --      clock_reset.reset
			scl_pad_io => scl_exp_export,                                              --       export_scl.export
			sda_pad_io => sda_exp_export,                                              --       export_sda.export
			wb_adr_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_opencores_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => i2c_opencores_0_interrupt_sender_irq                         -- interrupt_sender.irq
		);

	leds : component lms_orca_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_external_connection_export            -- external_connection.export
		);

	lms_ctr_gpio : component lms_orca_lms_ctr_gpio
		port map (
			clk        => clk_clk,                                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_lms_ctr_gpio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_lms_ctr_gpio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_lms_ctr_gpio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_lms_ctr_gpio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_lms_ctr_gpio_s1_readdata,        --                    .readdata
			out_port   => lms_ctr_gpio_external_connection_export            -- external_connection.export
		);

	oc_mem : component lms_orca_oc_mem
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_oc_mem_s1_address,    --     s1.address
			clken      => mm_interconnect_0_oc_mem_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_oc_mem_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_oc_mem_s1_write,      --       .write
			readdata   => mm_interconnect_0_oc_mem_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_oc_mem_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_oc_mem_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req      --       .reset_req
		);

	spi_1_dac : component lms_orca_spi_1_DAC
		port map (
			clk           => clk_clk,                                                      --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                     --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_1_dac_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_1_dac_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_1_dac_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_1_dac_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_1_dac_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_1_dac_spi_control_port_write_ports_inv, --                 .write_n
			irq           => spi_1_dac_irq_irq,                                            --              irq.irq
			MISO          => spi_1_dac_external_MISO,                                      --         external.export
			MOSI          => spi_1_dac_external_MOSI,                                      --                 .export
			SCLK          => spi_1_dac_external_SCLK,                                      --                 .export
			SS_n          => spi_1_dac_external_SS_n                                       --                 .export
		);

	spi_lms : component lms_orca_spi_lms
		port map (
			clk           => clk_clk,                                                    --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                   --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_lms_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_lms_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_lms_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_lms_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_lms_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_lms_spi_control_port_write_ports_inv, --                 .write_n
			irq           => spi_lms_irq_irq,                                            --              irq.irq
			MISO          => spi_lms_external_MISO,                                      --         external.export
			MOSI          => spi_lms_external_MOSI,                                      --                 .export
			SCLK          => spi_lms_external_SCLK,                                      --                 .export
			SS_n          => spi_lms_external_SS_n                                       --                 .export
		);

	switch : component lms_orca_switch
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_external_connection_export         -- external_connection.export
		);

	sysid_qsys_0 : component lms_orca_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	vectorblox_orca_0 : component Orca
		generic map (
			REGISTER_SIZE         => 32,
			AVALON_ENABLE         => 1,
			AXI_ENABLE            => 0,
			LVE_ENABLE            => 0,
			SCRATCHPAD_SIZE       => 1024,
			RESET_VECTOR          => 512,
			MULTIPLY_ENABLE       => 1,
			DIVIDE_ENABLE         => 0,
			SHIFTER_MAX_CYCLES    => 32,
			ENABLE_EXCEPTIONS     => 1,
			NUM_EXT_INTERRUPTS    => 1,
			ENABLE_EXT_INTERRUPTS => 1,
			COUNTER_LENGTH        => 64,
			BRANCH_PREDICTORS     => 1,
			PIPELINE_STAGES       => 4
		)
		port map (
			clk                           => clk_clk,                                     --             clock.clk
			scratchpad_clk                => clk_clk,                                     --    scratchpad_clk.clk
			reset                         => rst_controller_reset_out_reset,              --             reset.reset
			avm_data_address              => vectorblox_orca_0_data_address,              --              data.address
			avm_data_byteenable           => vectorblox_orca_0_data_byteenable,           --                  .byteenable
			avm_data_read                 => vectorblox_orca_0_data_read,                 --                  .read
			avm_data_readdata             => vectorblox_orca_0_data_readdata,             --                  .readdata
			avm_data_write                => vectorblox_orca_0_data_write,                --                  .write
			avm_data_writedata            => vectorblox_orca_0_data_writedata,            --                  .writedata
			avm_data_waitrequest          => vectorblox_orca_0_data_waitrequest,          --                  .waitrequest
			avm_data_readdatavalid        => vectorblox_orca_0_data_readdatavalid,        --                  .readdatavalid
			data_ARADDR                   => open,                                        --   axi_data_master.araddr
			data_ARBURST                  => open,                                        --                  .arburst
			data_ARCACHE                  => open,                                        --                  .arcache
			data_ARID                     => open,                                        --                  .arid
			data_ARLEN                    => open,                                        --                  .arlen
			data_ARLOCK                   => open,                                        --                  .arlock
			data_ARPROT                   => open,                                        --                  .arprot
			data_ARREADY                  => open,                                        --                  .arready
			data_ARSIZE                   => open,                                        --                  .arsize
			data_ARVALID                  => open,                                        --                  .arvalid
			data_AWADDR                   => open,                                        --                  .awaddr
			data_AWBURST                  => open,                                        --                  .awburst
			data_AWCACHE                  => open,                                        --                  .awcache
			data_AWID                     => open,                                        --                  .awid
			data_AWLEN                    => open,                                        --                  .awlen
			data_AWLOCK                   => open,                                        --                  .awlock
			data_AWPROT                   => open,                                        --                  .awprot
			data_AWREADY                  => open,                                        --                  .awready
			data_AWSIZE                   => open,                                        --                  .awsize
			data_AWVALID                  => open,                                        --                  .awvalid
			data_BID                      => open,                                        --                  .bid
			data_BREADY                   => open,                                        --                  .bready
			data_BRESP                    => open,                                        --                  .bresp
			data_BVALID                   => open,                                        --                  .bvalid
			data_RDATA                    => open,                                        --                  .rdata
			data_RID                      => open,                                        --                  .rid
			data_RLAST                    => open,                                        --                  .rlast
			data_RREADY                   => open,                                        --                  .rready
			data_RRESP                    => open,                                        --                  .rresp
			data_RVALID                   => open,                                        --                  .rvalid
			data_WDATA                    => open,                                        --                  .wdata
			data_WID                      => open,                                        --                  .wid
			data_WLAST                    => open,                                        --                  .wlast
			data_WREADY                   => open,                                        --                  .wready
			data_WSTRB                    => open,                                        --                  .wstrb
			data_WVALID                   => open,                                        --                  .wvalid
			instr_ARADDR                  => open,                                        --  axi_instr_master.araddr
			instr_ARBURST                 => open,                                        --                  .arburst
			instr_ARCACHE                 => open,                                        --                  .arcache
			instr_ARID                    => open,                                        --                  .arid
			instr_ARLEN                   => open,                                        --                  .arlen
			instr_ARLOCK                  => open,                                        --                  .arlock
			instr_ARPROT                  => open,                                        --                  .arprot
			instr_ARREADY                 => open,                                        --                  .arready
			instr_ARSIZE                  => open,                                        --                  .arsize
			instr_ARVALID                 => open,                                        --                  .arvalid
			instr_AWADDR                  => open,                                        --                  .awaddr
			instr_AWBURST                 => open,                                        --                  .awburst
			instr_AWCACHE                 => open,                                        --                  .awcache
			instr_AWID                    => open,                                        --                  .awid
			instr_AWLEN                   => open,                                        --                  .awlen
			instr_AWLOCK                  => open,                                        --                  .awlock
			instr_AWPROT                  => open,                                        --                  .awprot
			instr_AWREADY                 => open,                                        --                  .awready
			instr_AWSIZE                  => open,                                        --                  .awsize
			instr_AWVALID                 => open,                                        --                  .awvalid
			instr_BID                     => open,                                        --                  .bid
			instr_BREADY                  => open,                                        --                  .bready
			instr_BRESP                   => open,                                        --                  .bresp
			instr_BVALID                  => open,                                        --                  .bvalid
			instr_RDATA                   => open,                                        --                  .rdata
			instr_RID                     => open,                                        --                  .rid
			instr_RLAST                   => open,                                        --                  .rlast
			instr_RREADY                  => open,                                        --                  .rready
			instr_RRESP                   => open,                                        --                  .rresp
			instr_RVALID                  => open,                                        --                  .rvalid
			instr_WDATA                   => open,                                        --                  .wdata
			instr_WID                     => open,                                        --                  .wid
			instr_WLAST                   => open,                                        --                  .wlast
			instr_WREADY                  => open,                                        --                  .wready
			instr_WSTRB                   => open,                                        --                  .wstrb
			instr_WVALID                  => open,                                        --                  .wvalid
			avm_instruction_address       => vectorblox_orca_0_instruction_address,       --       instruction.address
			avm_instruction_read          => vectorblox_orca_0_instruction_read,          --                  .read
			avm_instruction_readdata      => vectorblox_orca_0_instruction_readdata,      --                  .readdata
			avm_instruction_waitrequest   => vectorblox_orca_0_instruction_waitrequest,   --                  .waitrequest
			avm_instruction_readdatavalid => vectorblox_orca_0_instruction_readdatavalid, --                  .readdatavalid
			global_interrupts             => vectorblox_orca_0_global_interrupts_export,  -- global_interrupts.export
			data_ADR_O                    => open,                                        --       (terminated)
			data_DAT_I                    => "00000000000000000000000000000000",          --       (terminated)
			data_DAT_O                    => open,                                        --       (terminated)
			data_WE_O                     => open,                                        --       (terminated)
			data_SEL_O                    => open,                                        --       (terminated)
			data_STB_O                    => open,                                        --       (terminated)
			data_ACK_I                    => '0',                                         --       (terminated)
			data_CYC_O                    => open,                                        --       (terminated)
			data_CTI_O                    => open,                                        --       (terminated)
			data_STALL_I                  => '0',                                         --       (terminated)
			instr_ADR_O                   => open,                                        --       (terminated)
			instr_DAT_I                   => "00000000000000000000000000000000",          --       (terminated)
			instr_STB_O                   => open,                                        --       (terminated)
			instr_ACK_I                   => '0',                                         --       (terminated)
			instr_CYC_O                   => open,                                        --       (terminated)
			instr_CTI_O                   => open,                                        --       (terminated)
			instr_STALL_I                 => '0'                                          --       (terminated)
		);

	mm_interconnect_0 : component lms_orca_mm_interconnect_0
		port map (
			clk_main_clk_clk                                    => clk_clk,                                                     --                                  clk_main_clk.clk
			vectorblox_orca_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- vectorblox_orca_0_reset_reset_bridge_in_reset.reset
			vectorblox_orca_0_data_address                      => vectorblox_orca_0_data_address,                              --                        vectorblox_orca_0_data.address
			vectorblox_orca_0_data_waitrequest                  => vectorblox_orca_0_data_waitrequest,                          --                                              .waitrequest
			vectorblox_orca_0_data_byteenable                   => vectorblox_orca_0_data_byteenable,                           --                                              .byteenable
			vectorblox_orca_0_data_read                         => vectorblox_orca_0_data_read,                                 --                                              .read
			vectorblox_orca_0_data_readdata                     => vectorblox_orca_0_data_readdata,                             --                                              .readdata
			vectorblox_orca_0_data_readdatavalid                => vectorblox_orca_0_data_readdatavalid,                        --                                              .readdatavalid
			vectorblox_orca_0_data_write                        => vectorblox_orca_0_data_write,                                --                                              .write
			vectorblox_orca_0_data_writedata                    => vectorblox_orca_0_data_writedata,                            --                                              .writedata
			vectorblox_orca_0_instruction_address               => vectorblox_orca_0_instruction_address,                       --                 vectorblox_orca_0_instruction.address
			vectorblox_orca_0_instruction_waitrequest           => vectorblox_orca_0_instruction_waitrequest,                   --                                              .waitrequest
			vectorblox_orca_0_instruction_read                  => vectorblox_orca_0_instruction_read,                          --                                              .read
			vectorblox_orca_0_instruction_readdata              => vectorblox_orca_0_instruction_readdata,                      --                                              .readdata
			vectorblox_orca_0_instruction_readdatavalid         => vectorblox_orca_0_instruction_readdatavalid,                 --                                              .readdatavalid
			Av_FIFO_Int_0_avalon_slave_0_address                => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address,      --                  Av_FIFO_Int_0_avalon_slave_0.address
			Av_FIFO_Int_0_avalon_slave_0_write                  => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write,        --                                              .write
			Av_FIFO_Int_0_avalon_slave_0_read                   => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read,         --                                              .read
			Av_FIFO_Int_0_avalon_slave_0_readdata               => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata,     --                                              .readdata
			Av_FIFO_Int_0_avalon_slave_0_writedata              => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata,    --                                              .writedata
			Av_FIFO_Int_0_avalon_slave_0_chipselect             => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect,   --                                              .chipselect
			controlled_reset_s1_address                         => mm_interconnect_0_controlled_reset_s1_address,               --                           controlled_reset_s1.address
			controlled_reset_s1_write                           => mm_interconnect_0_controlled_reset_s1_write,                 --                                              .write
			controlled_reset_s1_readdata                        => mm_interconnect_0_controlled_reset_s1_readdata,              --                                              .readdata
			controlled_reset_s1_writedata                       => mm_interconnect_0_controlled_reset_s1_writedata,             --                                              .writedata
			controlled_reset_s1_chipselect                      => mm_interconnect_0_controlled_reset_s1_chipselect,            --                                              .chipselect
			i2c_opencores_0_avalon_slave_0_address              => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --                i2c_opencores_0_avalon_slave_0.address
			i2c_opencores_0_avalon_slave_0_write                => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                                              .write
			i2c_opencores_0_avalon_slave_0_readdata             => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                                              .readdata
			i2c_opencores_0_avalon_slave_0_writedata            => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                                              .writedata
			i2c_opencores_0_avalon_slave_0_waitrequest          => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv,        --                                              .waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect           => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                                              .chipselect
			leds_s1_address                                     => mm_interconnect_0_leds_s1_address,                           --                                       leds_s1.address
			leds_s1_write                                       => mm_interconnect_0_leds_s1_write,                             --                                              .write
			leds_s1_readdata                                    => mm_interconnect_0_leds_s1_readdata,                          --                                              .readdata
			leds_s1_writedata                                   => mm_interconnect_0_leds_s1_writedata,                         --                                              .writedata
			leds_s1_chipselect                                  => mm_interconnect_0_leds_s1_chipselect,                        --                                              .chipselect
			lms_ctr_gpio_s1_address                             => mm_interconnect_0_lms_ctr_gpio_s1_address,                   --                               lms_ctr_gpio_s1.address
			lms_ctr_gpio_s1_write                               => mm_interconnect_0_lms_ctr_gpio_s1_write,                     --                                              .write
			lms_ctr_gpio_s1_readdata                            => mm_interconnect_0_lms_ctr_gpio_s1_readdata,                  --                                              .readdata
			lms_ctr_gpio_s1_writedata                           => mm_interconnect_0_lms_ctr_gpio_s1_writedata,                 --                                              .writedata
			lms_ctr_gpio_s1_chipselect                          => mm_interconnect_0_lms_ctr_gpio_s1_chipselect,                --                                              .chipselect
			oc_mem_s1_address                                   => mm_interconnect_0_oc_mem_s1_address,                         --                                     oc_mem_s1.address
			oc_mem_s1_write                                     => mm_interconnect_0_oc_mem_s1_write,                           --                                              .write
			oc_mem_s1_readdata                                  => mm_interconnect_0_oc_mem_s1_readdata,                        --                                              .readdata
			oc_mem_s1_writedata                                 => mm_interconnect_0_oc_mem_s1_writedata,                       --                                              .writedata
			oc_mem_s1_byteenable                                => mm_interconnect_0_oc_mem_s1_byteenable,                      --                                              .byteenable
			oc_mem_s1_chipselect                                => mm_interconnect_0_oc_mem_s1_chipselect,                      --                                              .chipselect
			oc_mem_s1_clken                                     => mm_interconnect_0_oc_mem_s1_clken,                           --                                              .clken
			spi_1_DAC_spi_control_port_address                  => mm_interconnect_0_spi_1_dac_spi_control_port_address,        --                    spi_1_DAC_spi_control_port.address
			spi_1_DAC_spi_control_port_write                    => mm_interconnect_0_spi_1_dac_spi_control_port_write,          --                                              .write
			spi_1_DAC_spi_control_port_read                     => mm_interconnect_0_spi_1_dac_spi_control_port_read,           --                                              .read
			spi_1_DAC_spi_control_port_readdata                 => mm_interconnect_0_spi_1_dac_spi_control_port_readdata,       --                                              .readdata
			spi_1_DAC_spi_control_port_writedata                => mm_interconnect_0_spi_1_dac_spi_control_port_writedata,      --                                              .writedata
			spi_1_DAC_spi_control_port_chipselect               => mm_interconnect_0_spi_1_dac_spi_control_port_chipselect,     --                                              .chipselect
			spi_lms_spi_control_port_address                    => mm_interconnect_0_spi_lms_spi_control_port_address,          --                      spi_lms_spi_control_port.address
			spi_lms_spi_control_port_write                      => mm_interconnect_0_spi_lms_spi_control_port_write,            --                                              .write
			spi_lms_spi_control_port_read                       => mm_interconnect_0_spi_lms_spi_control_port_read,             --                                              .read
			spi_lms_spi_control_port_readdata                   => mm_interconnect_0_spi_lms_spi_control_port_readdata,         --                                              .readdata
			spi_lms_spi_control_port_writedata                  => mm_interconnect_0_spi_lms_spi_control_port_writedata,        --                                              .writedata
			spi_lms_spi_control_port_chipselect                 => mm_interconnect_0_spi_lms_spi_control_port_chipselect,       --                                              .chipselect
			switch_s1_address                                   => mm_interconnect_0_switch_s1_address,                         --                                     switch_s1.address
			switch_s1_readdata                                  => mm_interconnect_0_switch_s1_readdata,                        --                                              .readdata
			sysid_qsys_0_control_slave_address                  => mm_interconnect_0_sysid_qsys_0_control_slave_address,        --                    sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                 => mm_interconnect_0_sysid_qsys_0_control_slave_readdata        --                                              .readdata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => in_reset_reset_n_ports_inv,         -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	in_reset_reset_n_ports_inv <= not in_reset_reset_n;

	mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv <= not i2c_opencores_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_lms_ctr_gpio_s1_write_ports_inv <= not mm_interconnect_0_lms_ctr_gpio_s1_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_controlled_reset_s1_write_ports_inv <= not mm_interconnect_0_controlled_reset_s1_write;

	mm_interconnect_0_spi_1_dac_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_1_dac_spi_control_port_read;

	mm_interconnect_0_spi_1_dac_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_1_dac_spi_control_port_write;

	mm_interconnect_0_spi_lms_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_lms_spi_control_port_read;

	mm_interconnect_0_spi_lms_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_lms_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of lms_orca
