
module clkctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
