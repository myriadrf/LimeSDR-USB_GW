@00000000
15000000
	 
